`timescale 1ns / 1ps

module kare_alici_4bit(
    input [3:0] a,
    output [7:0] f );
    
    assign f[0] = a[0];
    assign f[1] = ~a[0]&a[0];
    assign f[2] = (a[3]&a[2]&a[1]&(~a[0])) | (a[3]&(~a[2])&a[1]&(~a[0])) | ((~a[3])&a[2]&a[1]&(~a[0])) | ((~a[3])&(~a[2])&a[1]&(~a[0]));
    assign f[3] = (a[3]&a[2]&(~a[1])&a[0]) | (a[3]&(~a[2])&a[1]&a[0]) | ((~a[3])&a[2]&(~a[1])&a[0]) | ((~a[3])&(~a[2])&a[1]&a[0]);
    assign f[4] = (a[3]&a[2]&(~a[1])&(~a[0])) | (a[3]&(~a[2])&a[1]&a[0]) | (a[3]&(~a[2])&(~a[1])&a[0]) | ((~a[3])&a[2]&a[1]&a[0]) | ((~a[3])&a[2]&(~a[1])&a[0]) | ((~a[3])&a[2]&(~a[1])&(~a[0]));
    assign f[5] = (a[3]&a[2]&a[1]&a[0]) | (a[3]&a[2]&(~a[1])&a[0]) | (a[3]&(~a[2])&a[1]&a[0]) | (a[3]&(~a[2])&a[1]&(~a[0])) | ((~a[3])&a[2]&a[1]&a[0]) | ((~a[3])&a[2]&a[1]&(~a[0]));
    assign f[6] = (a[3]&a[2]&a[1]&a[0]) | (a[3]&a[2]&a[1]&(~a[0])) | (a[3]&(~a[2])&a[1]&a[0]) | (a[3]&(~a[2])&a[1]&(~a[0])) | (a[3]&(~a[2])&(~a[1])&a[0]) | (a[3]&(~a[2])&(~a[1])&(~a[0]));
    assign f[7] = (a[3]&a[2]&a[1]&a[0]) | (a[3]&a[2]&a[1]&(~a[0])) | (a[3]&a[2]&(~a[1])&a[0]) | (a[3]&a[2]&(~a[1])&(~a[0]));
    
endmodule
